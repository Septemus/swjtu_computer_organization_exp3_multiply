library verilog;
use verilog.vl_types.all;
entity keymodule_vlg_vec_tst is
end keymodule_vlg_vec_tst;
