library verilog;
use verilog.vl_types.all;
entity exp3_2_vlg_vec_tst is
end exp3_2_vlg_vec_tst;
